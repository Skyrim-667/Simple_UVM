`include "./verif/my_interface.sv"
`include "./coverage/coverage_collector.sv"
`include "./verif/transaction.sv"
`include "./verif/monitor_in.sv"
`include "./verif/monitor_out.sv"
`include "./verif/sequence.sv"
`include "./verif/sequencer.sv"
`include "./verif/vseqr.sv"
`include "./verif/vseq.sv"
`include "./verif/driver.sv"
`include "./verif/agent_in.sv"
`include "./verif/agent_out.sv"
`include "./verif/scb.sv"
`include "./verif/ref_model.sv"
`include "./verif/env.sv"
`include "./test_case/base_test.sv"
`include "./test_case/testcase_0.sv"


















